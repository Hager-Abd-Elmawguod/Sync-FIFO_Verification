package shared_pkg;
int error_count,correct_count;
event trigger;
endpackage